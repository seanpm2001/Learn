string S1 = "String"
